module cpu19 (
    input wire clk,
    input wire reset
);

//Program Counter
   reg[18:0] pc;
//pipeline registers
reg [18:0] instr_reg, alu_out_reg, memory_out_reg;
reg [18:0] reg_rs1, reg_rs2;
reg [18:0] reg_file_out1, regfile_rs2;
wire [18:0] alu_result;
wire alu_zero;
wire [4:0]opcode;
wire[3:0]rd, rs1, rs2;
wire [9:0] imm;
wire [13:0] addr;

wire fft_done;

    // Instantiate Control Unit
    control_unit CU (
        .instr(instr_reg),
        .opcode(opcode),
        .rd(rd),
        .rs1(rs1),
        .rs2(rs2),
        .imm(imm),
        .addr(addr)
    );

    // Instantiate Register File
    regfile RF (
        .clk(clk),
        .we(1'b0), // Placeholder, connect control logic
        .rd_addr(rd),
        .rs1_addr(rs1),
        .rs2_addr(rs2),
        .wd(alu_result),
        .rs1(regfile_out1),
        .rs2(regfile_out2)
    );

    // Instantiate ALU
    alu ALU (
        .opcode(opcode),
        .a(regfile_out1),
        .b(regfile_out2),
        .result(alu_result),
        .zero(alu_zero)
    );

    // Instantiate FFT Accelerator
    fft_accel FFTU (
        .clk(clk),
        .start(1'b0), // Placeholder, connect control logic
        .addr_in(regfile_out2),
        .addr_out(regfile_out1),
        .done(fft_done)
    );

    // Instantiate Memory Interface
    wire [18:0] mem_data;
    wire [18:0] mem_out;
    mem_interface MEM (
        .clk(clk),
        .we(1'b0), // Placeholder, connect control logic
        .addr(alu_result),
        .data(mem_data),
        .mem_out(mem_out),
        .mem_in(regfile_out2)
    );

    // Instruction Fetch (placeholder)
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            pc <= 19'b0;
        end else begin
            // Fetch instruction from memory (placeholder)
            instr_reg <= mem_out;
            // Update PC (placeholder)
            pc <= pc + 1;
        end
    end
endmodule 
